library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity game_text is

	port (	draw_clk 	: in std_logic;

			win			: in std_logic;
			lose		: in std_logic;

			draw_x		: in integer range 0 to 319;
			draw_y		: in integer range 0 to 239;
			pixel		: out std_logic);

end game_text;

architecture behavioral of game_text is

	type sprite_t is array (9 downto 0) of std_logic_vector (75 downto 0);

	constant sprite_a : sprite_t := ("0000011000011000011110000110000110000000000110000110011111111001110001100000",
									 "0000011000011000111111000110000110000000000110000110011111111001110001100000",
									 "0000011000011001100001100110000110000000000110000110000011000001101001100000",
									 "0000011000011001100001100110000110000000000110000110000011000001101001100000",
									 "0000011000011001100001100110000110000000000110110110000011000001100101100000",
									 "0000001100110001100001100110000110000000000110110110000011000001100101100000",
									 "0000000111100001100001100110000110000000000110110110000011000001100011100000",
									 "0000000011000001100001100110000110000000000110110110000011000001100011100000",
									 "0000000011000000111111000011111100000000000011111100011111111001100001100000",
									 "0000000011000000011110000001111000000000000011001100011111111001100001100000");

	constant sprite_b : sprite_t := ("1100001100001111000011000011000000000011000000000011110000001111110001111111",
									 "1100001100011111100011000011000000000011000000000111111000011111110011111111",
									 "1100001100110000110011000011000000000011000000001100001100110000000011000000",
									 "1100001100110000110011000011000000000011000000001100001100110000000011000000",
									 "1100001100110000110011000011000000000011000000001100001100011111000001111000",
									 "0110011000110000110011000011000000000011000000001100001100001111100001111000",
									 "0011110000110000110011000011000000000011000000001100001100000000110011000000",
									 "0001100000110000110011000011000000000011000000001100001100000000110011000000",
									 "0001100000011111100001111110000000000011111111000111111000111111100011111111",
									 "0001100000001111000000111100000000000011111111000011110000111111000001111111");

	constant cx : integer := 122;
	constant cy : integer := 115;

	signal rx	: integer range -1 to 76;
	signal ry	: integer range -1 to 10;

begin

	--------------------------------------------------------------------------------------------------------------------
	-- DRAW

	rx <= (draw_x - cx) when ((draw_x >= cx) and (draw_x <= (cx + 75))) else -1;
	ry <= (draw_y - cy) when ((draw_y >= cy) and (draw_y <= (cy + 9))) else -1;

	draw_p : process (draw_clk)
	begin
		if rising_edge(draw_clk) then
			if ((rx = -1) or (ry = -1)) then
				pixel <= '0';
			elsif (win = '1') then
				pixel <= sprite_a (9 - ry) (75 - rx);
			elsif (lose = '1') then
				pixel <= sprite_b (9 - ry) (75 - rx);
			else
				pixel <= '0';
			end if;
		end if;
	end process;

end behavioral;